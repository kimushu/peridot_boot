// ngs_boot_core.v

// Generated using ACDS version 16.1 203

`timescale 1 ps / 1 ps
module ngs_boot_core (
		input  wire        clk_100m_clk,           // clk_100m.clk
		input  wire        clk_25m_clk,            //  clk_25m.clk
		output wire        epcs_cso_n,             //     epcs.cso_n
		output wire        epcs_dclk,              //         .dclk
		output wire        epcs_asdo,              //         .asdo
		input  wire        epcs_data0,             //         .data0
		inout  wire [29:0] gpio_export,            //     gpio.export
		input  wire        hostuart_rxd,           // hostuart.rxd
		output wire        hostuart_txd,           //         .txd
		input  wire        mreset_mreset_n,        //   mreset.mreset_n
		input  wire        nios2_cpu_resetrequest, //    nios2.cpu_resetrequest
		output wire        nios2_cpu_resettaken,   //         .cpu_resettaken
		input  wire        reset_reset_n,          //    reset.reset_n
		output wire [11:0] sdr_addr,               //      sdr.addr
		output wire [1:0]  sdr_ba,                 //         .ba
		output wire        sdr_cas_n,              //         .cas_n
		output wire        sdr_cke,                //         .cke
		output wire        sdr_cs_n,               //         .cs_n
		inout  wire [15:0] sdr_dq,                 //         .dq
		output wire [1:0]  sdr_dqm,                //         .dqm
		output wire        sdr_ras_n,              //         .ras_n
		output wire        sdr_we_n,               //         .we_n
		output wire        swi_cpu_resetrequest,   //      swi.cpu_resetrequest
		output wire [3:0]  swi_led                 //         .led
	);

	wire  [31:0] nios2_fast_data_master_readdata;                           // mm_interconnect_0:nios2_fast_data_master_readdata -> nios2_fast:d_readdata
	wire         nios2_fast_data_master_waitrequest;                        // mm_interconnect_0:nios2_fast_data_master_waitrequest -> nios2_fast:d_waitrequest
	wire         nios2_fast_data_master_debugaccess;                        // nios2_fast:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_fast_data_master_debugaccess
	wire  [28:0] nios2_fast_data_master_address;                            // nios2_fast:d_address -> mm_interconnect_0:nios2_fast_data_master_address
	wire   [3:0] nios2_fast_data_master_byteenable;                         // nios2_fast:d_byteenable -> mm_interconnect_0:nios2_fast_data_master_byteenable
	wire         nios2_fast_data_master_read;                               // nios2_fast:d_read -> mm_interconnect_0:nios2_fast_data_master_read
	wire         nios2_fast_data_master_readdatavalid;                      // mm_interconnect_0:nios2_fast_data_master_readdatavalid -> nios2_fast:d_readdatavalid
	wire         nios2_fast_data_master_write;                              // nios2_fast:d_write -> mm_interconnect_0:nios2_fast_data_master_write
	wire  [31:0] nios2_fast_data_master_writedata;                          // nios2_fast:d_writedata -> mm_interconnect_0:nios2_fast_data_master_writedata
	wire  [31:0] peridot_hostbridge_m1_readdata;                            // mm_interconnect_0:peridot_hostbridge_m1_readdata -> peridot_hostbridge:avm_m1_readdata
	wire         peridot_hostbridge_m1_waitrequest;                         // mm_interconnect_0:peridot_hostbridge_m1_waitrequest -> peridot_hostbridge:avm_m1_waitrequest
	wire  [31:0] peridot_hostbridge_m1_address;                             // peridot_hostbridge:avm_m1_address -> mm_interconnect_0:peridot_hostbridge_m1_address
	wire         peridot_hostbridge_m1_read;                                // peridot_hostbridge:avm_m1_read -> mm_interconnect_0:peridot_hostbridge_m1_read
	wire   [3:0] peridot_hostbridge_m1_byteenable;                          // peridot_hostbridge:avm_m1_byteenable -> mm_interconnect_0:peridot_hostbridge_m1_byteenable
	wire         peridot_hostbridge_m1_readdatavalid;                       // mm_interconnect_0:peridot_hostbridge_m1_readdatavalid -> peridot_hostbridge:avm_m1_readdatavalid
	wire         peridot_hostbridge_m1_write;                               // peridot_hostbridge:avm_m1_write -> mm_interconnect_0:peridot_hostbridge_m1_write
	wire  [31:0] peridot_hostbridge_m1_writedata;                           // peridot_hostbridge:avm_m1_writedata -> mm_interconnect_0:peridot_hostbridge_m1_writedata
	wire  [31:0] nios2_fast_instruction_master_readdata;                    // mm_interconnect_0:nios2_fast_instruction_master_readdata -> nios2_fast:i_readdata
	wire         nios2_fast_instruction_master_waitrequest;                 // mm_interconnect_0:nios2_fast_instruction_master_waitrequest -> nios2_fast:i_waitrequest
	wire  [27:0] nios2_fast_instruction_master_address;                     // nios2_fast:i_address -> mm_interconnect_0:nios2_fast_instruction_master_address
	wire         nios2_fast_instruction_master_read;                        // nios2_fast:i_read -> mm_interconnect_0:nios2_fast_instruction_master_read
	wire         nios2_fast_instruction_master_readdatavalid;               // mm_interconnect_0:nios2_fast_instruction_master_readdatavalid -> nios2_fast:i_readdatavalid
	wire  [31:0] mm_interconnect_0_ufm_data_readdata;                       // ufm:avmm_data_readdata -> mm_interconnect_0:ufm_data_readdata
	wire         mm_interconnect_0_ufm_data_waitrequest;                    // ufm:avmm_data_waitrequest -> mm_interconnect_0:ufm_data_waitrequest
	wire  [15:0] mm_interconnect_0_ufm_data_address;                        // mm_interconnect_0:ufm_data_address -> ufm:avmm_data_addr
	wire         mm_interconnect_0_ufm_data_read;                           // mm_interconnect_0:ufm_data_read -> ufm:avmm_data_read
	wire         mm_interconnect_0_ufm_data_readdatavalid;                  // ufm:avmm_data_readdatavalid -> mm_interconnect_0:ufm_data_readdatavalid
	wire         mm_interconnect_0_ufm_data_write;                          // mm_interconnect_0:ufm_data_write -> ufm:avmm_data_write
	wire  [31:0] mm_interconnect_0_ufm_data_writedata;                      // mm_interconnect_0:ufm_data_writedata -> ufm:avmm_data_writedata
	wire   [1:0] mm_interconnect_0_ufm_data_burstcount;                     // mm_interconnect_0:ufm_data_burstcount -> ufm:avmm_data_burstcount
	wire  [31:0] mm_interconnect_0_nios2_fast_debug_mem_slave_readdata;     // nios2_fast:debug_mem_slave_readdata -> mm_interconnect_0:nios2_fast_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_fast_debug_mem_slave_waitrequest;  // nios2_fast:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_fast_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_fast_debug_mem_slave_debugaccess;  // mm_interconnect_0:nios2_fast_debug_mem_slave_debugaccess -> nios2_fast:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_fast_debug_mem_slave_address;      // mm_interconnect_0:nios2_fast_debug_mem_slave_address -> nios2_fast:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_fast_debug_mem_slave_read;         // mm_interconnect_0:nios2_fast_debug_mem_slave_read -> nios2_fast:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_fast_debug_mem_slave_byteenable;   // mm_interconnect_0:nios2_fast_debug_mem_slave_byteenable -> nios2_fast:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_fast_debug_mem_slave_write;        // mm_interconnect_0:nios2_fast_debug_mem_slave_write -> nios2_fast:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_fast_debug_mem_slave_writedata;    // mm_interconnect_0:nios2_fast_debug_mem_slave_writedata -> nios2_fast:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_peripheral_bridge_s0_readdata;           // peripheral_bridge:s0_readdata -> mm_interconnect_0:peripheral_bridge_s0_readdata
	wire         mm_interconnect_0_peripheral_bridge_s0_waitrequest;        // peripheral_bridge:s0_waitrequest -> mm_interconnect_0:peripheral_bridge_s0_waitrequest
	wire         mm_interconnect_0_peripheral_bridge_s0_debugaccess;        // mm_interconnect_0:peripheral_bridge_s0_debugaccess -> peripheral_bridge:s0_debugaccess
	wire  [15:0] mm_interconnect_0_peripheral_bridge_s0_address;            // mm_interconnect_0:peripheral_bridge_s0_address -> peripheral_bridge:s0_address
	wire         mm_interconnect_0_peripheral_bridge_s0_read;               // mm_interconnect_0:peripheral_bridge_s0_read -> peripheral_bridge:s0_read
	wire   [3:0] mm_interconnect_0_peripheral_bridge_s0_byteenable;         // mm_interconnect_0:peripheral_bridge_s0_byteenable -> peripheral_bridge:s0_byteenable
	wire         mm_interconnect_0_peripheral_bridge_s0_readdatavalid;      // peripheral_bridge:s0_readdatavalid -> mm_interconnect_0:peripheral_bridge_s0_readdatavalid
	wire         mm_interconnect_0_peripheral_bridge_s0_write;              // mm_interconnect_0:peripheral_bridge_s0_write -> peripheral_bridge:s0_write
	wire  [31:0] mm_interconnect_0_peripheral_bridge_s0_writedata;          // mm_interconnect_0:peripheral_bridge_s0_writedata -> peripheral_bridge:s0_writedata
	wire   [0:0] mm_interconnect_0_peripheral_bridge_s0_burstcount;         // mm_interconnect_0:peripheral_bridge_s0_burstcount -> peripheral_bridge:s0_burstcount
	wire         mm_interconnect_0_sdram_s1_chipselect;                     // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;                       // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                    // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [21:0] mm_interconnect_0_sdram_s1_address;                        // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                           // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;                     // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                  // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                          // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;                      // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire         peripheral_bridge_m0_waitrequest;                          // mm_interconnect_1:peripheral_bridge_m0_waitrequest -> peripheral_bridge:m0_waitrequest
	wire  [31:0] peripheral_bridge_m0_readdata;                             // mm_interconnect_1:peripheral_bridge_m0_readdata -> peripheral_bridge:m0_readdata
	wire         peripheral_bridge_m0_debugaccess;                          // peripheral_bridge:m0_debugaccess -> mm_interconnect_1:peripheral_bridge_m0_debugaccess
	wire  [15:0] peripheral_bridge_m0_address;                              // peripheral_bridge:m0_address -> mm_interconnect_1:peripheral_bridge_m0_address
	wire         peripheral_bridge_m0_read;                                 // peripheral_bridge:m0_read -> mm_interconnect_1:peripheral_bridge_m0_read
	wire   [3:0] peripheral_bridge_m0_byteenable;                           // peripheral_bridge:m0_byteenable -> mm_interconnect_1:peripheral_bridge_m0_byteenable
	wire         peripheral_bridge_m0_readdatavalid;                        // mm_interconnect_1:peripheral_bridge_m0_readdatavalid -> peripheral_bridge:m0_readdatavalid
	wire  [31:0] peripheral_bridge_m0_writedata;                            // peripheral_bridge:m0_writedata -> mm_interconnect_1:peripheral_bridge_m0_writedata
	wire         peripheral_bridge_m0_write;                                // peripheral_bridge:m0_write -> mm_interconnect_1:peripheral_bridge_m0_write
	wire   [0:0] peripheral_bridge_m0_burstcount;                           // peripheral_bridge:m0_burstcount -> mm_interconnect_1:peripheral_bridge_m0_burstcount
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_1:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata;    // jtag_uart:av_readdata -> mm_interconnect_1:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest; // jtag_uart:av_waitrequest -> mm_interconnect_1:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_1:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_1:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_1:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_1:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_1_ufm_csr_readdata;                        // ufm:avmm_csr_readdata -> mm_interconnect_1:ufm_csr_readdata
	wire   [0:0] mm_interconnect_1_ufm_csr_address;                         // mm_interconnect_1:ufm_csr_address -> ufm:avmm_csr_addr
	wire         mm_interconnect_1_ufm_csr_read;                            // mm_interconnect_1:ufm_csr_read -> ufm:avmm_csr_read
	wire         mm_interconnect_1_ufm_csr_write;                           // mm_interconnect_1:ufm_csr_write -> ufm:avmm_csr_write
	wire  [31:0] mm_interconnect_1_ufm_csr_writedata;                       // mm_interconnect_1:ufm_csr_writedata -> ufm:avmm_csr_writedata
	wire         mm_interconnect_1_systimer_s1_chipselect;                  // mm_interconnect_1:systimer_s1_chipselect -> systimer:chipselect
	wire  [15:0] mm_interconnect_1_systimer_s1_readdata;                    // systimer:readdata -> mm_interconnect_1:systimer_s1_readdata
	wire   [2:0] mm_interconnect_1_systimer_s1_address;                     // mm_interconnect_1:systimer_s1_address -> systimer:address
	wire         mm_interconnect_1_systimer_s1_write;                       // mm_interconnect_1:systimer_s1_write -> systimer:write_n
	wire  [15:0] mm_interconnect_1_systimer_s1_writedata;                   // mm_interconnect_1:systimer_s1_writedata -> systimer:writedata
	wire  [31:0] mm_interconnect_1_peridot_hostbridge_s1_readdata;          // peridot_hostbridge:avs_s1_readdata -> mm_interconnect_1:peridot_hostbridge_s1_readdata
	wire   [2:0] mm_interconnect_1_peridot_hostbridge_s1_address;           // mm_interconnect_1:peridot_hostbridge_s1_address -> peridot_hostbridge:avs_s1_address
	wire         mm_interconnect_1_peridot_hostbridge_s1_read;              // mm_interconnect_1:peridot_hostbridge_s1_read -> peridot_hostbridge:avs_s1_read
	wire         mm_interconnect_1_peridot_hostbridge_s1_write;             // mm_interconnect_1:peridot_hostbridge_s1_write -> peridot_hostbridge:avs_s1_write
	wire  [31:0] mm_interconnect_1_peridot_hostbridge_s1_writedata;         // mm_interconnect_1:peridot_hostbridge_s1_writedata -> peridot_hostbridge:avs_s1_writedata
	wire         mm_interconnect_1_gpio_s1_chipselect;                      // mm_interconnect_1:gpio_s1_chipselect -> gpio:chipselect
	wire  [31:0] mm_interconnect_1_gpio_s1_readdata;                        // gpio:readdata -> mm_interconnect_1:gpio_s1_readdata
	wire   [2:0] mm_interconnect_1_gpio_s1_address;                         // mm_interconnect_1:gpio_s1_address -> gpio:address
	wire         mm_interconnect_1_gpio_s1_write;                           // mm_interconnect_1:gpio_s1_write -> gpio:write_n
	wire  [31:0] mm_interconnect_1_gpio_s1_writedata;                       // mm_interconnect_1:gpio_s1_writedata -> gpio:writedata
	wire         irq_mapper_receiver0_irq;                                  // peridot_hostbridge:ins_avsirq_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver2_irq;                                  // jtag_uart:av_irq -> irq_mapper:receiver2_irq
	wire  [31:0] nios2_fast_irq_irq;                                        // irq_mapper:sender_irq -> nios2_fast:irq
	wire         irq_mapper_receiver1_irq;                                  // irq_synchronizer:sender_irq -> irq_mapper:receiver1_irq
	wire   [0:0] irq_synchronizer_receiver_irq;                             // systimer:irq -> irq_synchronizer:receiver_irq
	wire         irq_mapper_receiver3_irq;                                  // irq_synchronizer_001:sender_irq -> irq_mapper:receiver3_irq
	wire   [0:0] irq_synchronizer_001_receiver_irq;                         // gpio:irq -> irq_synchronizer_001:receiver_irq
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [gpio:reset_n, irq_synchronizer:receiver_reset, irq_synchronizer_001:receiver_reset, mm_interconnect_0:peripheral_bridge_reset_reset_bridge_in_reset_reset, mm_interconnect_1:peripheral_bridge_reset_reset_bridge_in_reset_reset, peridot_hostbridge:csi_avsclock_reset, peripheral_bridge:reset, systimer:reset_n]
	wire         rst_controller_001_reset_out_reset;                        // rst_controller_001:reset_out -> [jtag_uart:rst_n, mm_interconnect_1:jtag_uart_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_002_reset_out_reset;                        // rst_controller_002:reset_out -> [irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, mm_interconnect_0:nios2_fast_reset_reset_bridge_in_reset_reset, mm_interconnect_1:ufm_nreset_reset_bridge_in_reset_reset, nios2_fast:reset_n, peridot_hostbridge:csi_avmclock_reset, rst_translator:in_reset, sdram:reset_n, ufm:reset_n]
	wire         rst_controller_002_reset_out_reset_req;                    // rst_controller_002:reset_req -> [nios2_fast:reset_req, rst_translator:reset_req_in]

	ngs_boot_core_gpio gpio (
		.clk        (clk_25m_clk),                          //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_1_gpio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_gpio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_gpio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_gpio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_gpio_s1_readdata),   //                    .readdata
		.bidir_port (gpio_export),                          // external_connection.export
		.irq        (irq_synchronizer_001_receiver_irq)     //                 irq.irq
	);

	ngs_boot_core_jtag_uart jtag_uart (
		.clk            (clk_100m_clk),                                              //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_1_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_1_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_1_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver2_irq)                                   //               irq.irq
	);

	ngs_boot_core_nios2_fast nios2_fast (
		.clk                                 (clk_100m_clk),                                             //                       clk.clk
		.reset_n                             (~rst_controller_002_reset_out_reset),                      //                     reset.reset_n
		.reset_req                           (rst_controller_002_reset_out_reset_req),                   //                          .reset_req
		.d_address                           (nios2_fast_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_fast_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_fast_data_master_read),                              //                          .read
		.d_readdata                          (nios2_fast_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_fast_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_fast_data_master_write),                             //                          .write
		.d_writedata                         (nios2_fast_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (nios2_fast_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (nios2_fast_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_fast_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_fast_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_fast_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_fast_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (nios2_fast_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios2_fast_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                         //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_fast_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_fast_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_fast_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_fast_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_fast_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_fast_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_fast_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_fast_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       (),                                                         // custom_instruction_master.readra
		.cpu_resetrequest                    (nios2_cpu_resetrequest),                                   //  cpu_resetrequest_conduit.cpu_resetrequest
		.cpu_resettaken                      (nios2_cpu_resettaken)                                      //                          .cpu_resettaken
	);

	peridot_hostbridge #(
		.DEVICE_FAMILY        ("MAX 10"),
		.AVM_CLOCKFREQ        (100000000),
		.AVS_CLOCKFREQ        (25000000),
		.RECONFIG_FEATURE     ("DISABLE"),
		.INSTANCE_ALTDUALBOOT ("ENABLE"),
		.CHIPUID_FEATURE      ("ENABLE"),
		.HOSTINTERFACE_TYPE   ("UART"),
		.HOSTUART_BAUDRATE    (115200),
		.HOSTUART_INFIFODEPTH (6),
		.PERIDOT_GENCODE      (88),
		.RECONF_DELAY_CYCLE   (5000000),
		.CONFIG_CYCLE         (9),
		.RESET_TIMER_CYCLE    (13),
		.SWI_EPCSBOOT_FEATURE ("ENABLE"),
		.SWI_UIDREAD_FEATURE  ("ENABLE"),
		.SWI_MESSAGE_FEATURE  ("ENABLE"),
		.SWI_CLASSID          (32'b01110010101010010000000000000000),
		.SWI_TIMECODE         (1489088162),
		.SWI_CPURESET_KEY     (16'b1101111010101101),
		.SWI_CPURESET_INIT    (1)
	) peridot_hostbridge (
		.csi_avmclock_clk     (clk_100m_clk),                                      //  avmclock.clk
		.csi_avmclock_reset   (rst_controller_002_reset_out_reset),                //  avmreset.reset
		.avm_m1_address       (peridot_hostbridge_m1_address),                     //        m1.address
		.avm_m1_readdata      (peridot_hostbridge_m1_readdata),                    //          .readdata
		.avm_m1_read          (peridot_hostbridge_m1_read),                        //          .read
		.avm_m1_write         (peridot_hostbridge_m1_write),                       //          .write
		.avm_m1_byteenable    (peridot_hostbridge_m1_byteenable),                  //          .byteenable
		.avm_m1_writedata     (peridot_hostbridge_m1_writedata),                   //          .writedata
		.avm_m1_waitrequest   (peridot_hostbridge_m1_waitrequest),                 //          .waitrequest
		.avm_m1_readdatavalid (peridot_hostbridge_m1_readdatavalid),               //          .readdatavalid
		.csi_avsclock_clk     (clk_25m_clk),                                       //  avsclock.clk
		.csi_avsclock_reset   (rst_controller_reset_out_reset),                    //  avsreset.reset
		.avs_s1_address       (mm_interconnect_1_peridot_hostbridge_s1_address),   //        s1.address
		.avs_s1_read          (mm_interconnect_1_peridot_hostbridge_s1_read),      //          .read
		.avs_s1_readdata      (mm_interconnect_1_peridot_hostbridge_s1_readdata),  //          .readdata
		.avs_s1_write         (mm_interconnect_1_peridot_hostbridge_s1_write),     //          .write
		.avs_s1_writedata     (mm_interconnect_1_peridot_hostbridge_s1_writedata), //          .writedata
		.ins_avsirq_irq       (irq_mapper_receiver0_irq),                          //    avsirq.irq
		.rso_busreset_reset   (),                                                  //  busreset.reset
		.coe_mreset_n         (mreset_mreset_n),                                   // corereset.mreset_n
		.coe_rxd              (hostuart_rxd),                                      //  hostuart.rxd
		.coe_txd              (hostuart_txd),                                      //          .txd
		.coe_cpureset         (swi_cpu_resetrequest),                              //       swi.cpu_resetrequest
		.coe_led              (swi_led),                                           //          .led
		.coe_cso_n            (epcs_cso_n),                                        //  swi_epcs.cso_n
		.coe_dclk             (epcs_dclk),                                         //          .dclk
		.coe_asdo             (epcs_asdo),                                         //          .asdo
		.coe_data0            (epcs_data0),                                        //          .data0
		.coe_ft_d             (),                                                  // (terminated)
		.coe_ft_rd_n          (),                                                  // (terminated)
		.coe_ft_wr            (),                                                  // (terminated)
		.coe_ft_rxf_n         (1'b0),                                              // (terminated)
		.coe_ft_txe_n         (1'b0),                                              // (terminated)
		.coe_ft_siwu_n        ()                                                   // (terminated)
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (16),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) peripheral_bridge (
		.clk              (clk_25m_clk),                                          //   clk.clk
		.reset            (rst_controller_reset_out_reset),                       // reset.reset
		.s0_waitrequest   (mm_interconnect_0_peripheral_bridge_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_0_peripheral_bridge_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_0_peripheral_bridge_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_0_peripheral_bridge_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_0_peripheral_bridge_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_0_peripheral_bridge_s0_address),       //      .address
		.s0_write         (mm_interconnect_0_peripheral_bridge_s0_write),         //      .write
		.s0_read          (mm_interconnect_0_peripheral_bridge_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_0_peripheral_bridge_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_0_peripheral_bridge_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (peripheral_bridge_m0_waitrequest),                     //    m0.waitrequest
		.m0_readdata      (peripheral_bridge_m0_readdata),                        //      .readdata
		.m0_readdatavalid (peripheral_bridge_m0_readdatavalid),                   //      .readdatavalid
		.m0_burstcount    (peripheral_bridge_m0_burstcount),                      //      .burstcount
		.m0_writedata     (peripheral_bridge_m0_writedata),                       //      .writedata
		.m0_address       (peripheral_bridge_m0_address),                         //      .address
		.m0_write         (peripheral_bridge_m0_write),                           //      .write
		.m0_read          (peripheral_bridge_m0_read),                            //      .read
		.m0_byteenable    (peripheral_bridge_m0_byteenable),                      //      .byteenable
		.m0_debugaccess   (peripheral_bridge_m0_debugaccess),                     //      .debugaccess
		.s0_response      (),                                                     // (terminated)
		.m0_response      (2'b00)                                                 // (terminated)
	);

	ngs_boot_core_sdram sdram (
		.clk            (clk_100m_clk),                             //   clk.clk
		.reset_n        (~rst_controller_002_reset_out_reset),      // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdr_addr),                                 //  wire.export
		.zs_ba          (sdr_ba),                                   //      .export
		.zs_cas_n       (sdr_cas_n),                                //      .export
		.zs_cke         (sdr_cke),                                  //      .export
		.zs_cs_n        (sdr_cs_n),                                 //      .export
		.zs_dq          (sdr_dq),                                   //      .export
		.zs_dqm         (sdr_dqm),                                  //      .export
		.zs_ras_n       (sdr_ras_n),                                //      .export
		.zs_we_n        (sdr_we_n)                                  //      .export
	);

	ngs_boot_core_systimer systimer (
		.clk        (clk_25m_clk),                              //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          // reset.reset_n
		.address    (mm_interconnect_1_systimer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_1_systimer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_1_systimer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_1_systimer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_1_systimer_s1_write),     //      .write_n
		.irq        (irq_synchronizer_receiver_irq)             //   irq.irq
	);

	altera_onchip_flash #(
		.INIT_FILENAME                       (""),
		.INIT_FILENAME_SIM                   (""),
		.DEVICE_FAMILY                       ("MAX 10"),
		.PART_NAME                           ("10M08SAE144C8G"),
		.DEVICE_ID                           ("08"),
		.SECTOR1_START_ADDR                  (0),
		.SECTOR1_END_ADDR                    (4095),
		.SECTOR2_START_ADDR                  (4096),
		.SECTOR2_END_ADDR                    (8191),
		.SECTOR3_START_ADDR                  (8192),
		.SECTOR3_END_ADDR                    (29183),
		.SECTOR4_START_ADDR                  (29184),
		.SECTOR4_END_ADDR                    (44031),
		.SECTOR5_START_ADDR                  (0),
		.SECTOR5_END_ADDR                    (0),
		.MIN_VALID_ADDR                      (0),
		.MAX_VALID_ADDR                      (44031),
		.MIN_UFM_VALID_ADDR                  (0),
		.MAX_UFM_VALID_ADDR                  (8191),
		.SECTOR1_MAP                         (1),
		.SECTOR2_MAP                         (2),
		.SECTOR3_MAP                         (3),
		.SECTOR4_MAP                         (4),
		.SECTOR5_MAP                         (0),
		.ADDR_RANGE1_END_ADDR                (44031),
		.ADDR_RANGE1_OFFSET                  (512),
		.ADDR_RANGE2_OFFSET                  (0),
		.AVMM_DATA_ADDR_WIDTH                (16),
		.AVMM_DATA_DATA_WIDTH                (32),
		.AVMM_DATA_BURSTCOUNT_WIDTH          (2),
		.SECTOR_READ_PROTECTION_MODE         (16),
		.FLASH_SEQ_READ_DATA_COUNT           (2),
		.FLASH_ADDR_ALIGNMENT_BITS           (1),
		.FLASH_READ_CYCLE_MAX_INDEX          (4),
		.FLASH_RESET_CYCLE_MAX_INDEX         (25),
		.FLASH_BUSY_TIMEOUT_CYCLE_MAX_INDEX  (120),
		.FLASH_ERASE_TIMEOUT_CYCLE_MAX_INDEX (35000000),
		.FLASH_WRITE_TIMEOUT_CYCLE_MAX_INDEX (30500),
		.PARALLEL_MODE                       (1),
		.READ_AND_WRITE_MODE                 (1),
		.WRAPPING_BURST_MODE                 (0),
		.IS_DUAL_BOOT                        ("True"),
		.IS_ERAM_SKIP                        ("True"),
		.IS_COMPRESSED_IMAGE                 ("True")
	) ufm (
		.clock                   (clk_100m_clk),                             //    clk.clk
		.reset_n                 (~rst_controller_002_reset_out_reset),      // nreset.reset_n
		.avmm_data_addr          (mm_interconnect_0_ufm_data_address),       //   data.address
		.avmm_data_read          (mm_interconnect_0_ufm_data_read),          //       .read
		.avmm_data_writedata     (mm_interconnect_0_ufm_data_writedata),     //       .writedata
		.avmm_data_write         (mm_interconnect_0_ufm_data_write),         //       .write
		.avmm_data_readdata      (mm_interconnect_0_ufm_data_readdata),      //       .readdata
		.avmm_data_waitrequest   (mm_interconnect_0_ufm_data_waitrequest),   //       .waitrequest
		.avmm_data_readdatavalid (mm_interconnect_0_ufm_data_readdatavalid), //       .readdatavalid
		.avmm_data_burstcount    (mm_interconnect_0_ufm_data_burstcount),    //       .burstcount
		.avmm_csr_addr           (mm_interconnect_1_ufm_csr_address),        //    csr.address
		.avmm_csr_read           (mm_interconnect_1_ufm_csr_read),           //       .read
		.avmm_csr_writedata      (mm_interconnect_1_ufm_csr_writedata),      //       .writedata
		.avmm_csr_write          (mm_interconnect_1_ufm_csr_write),          //       .write
		.avmm_csr_readdata       (mm_interconnect_1_ufm_csr_readdata)        //       .readdata
	);

	ngs_boot_core_mm_interconnect_0 mm_interconnect_0 (
		.core_clk_clk_clk                                    (clk_100m_clk),                                             //                                  core_clk_clk.clk
		.peri_clk_clk_clk                                    (clk_25m_clk),                                              //                                  peri_clk_clk.clk
		.nios2_fast_reset_reset_bridge_in_reset_reset        (rst_controller_002_reset_out_reset),                       //        nios2_fast_reset_reset_bridge_in_reset.reset
		.peripheral_bridge_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                           // peripheral_bridge_reset_reset_bridge_in_reset.reset
		.nios2_fast_data_master_address                      (nios2_fast_data_master_address),                           //                        nios2_fast_data_master.address
		.nios2_fast_data_master_waitrequest                  (nios2_fast_data_master_waitrequest),                       //                                              .waitrequest
		.nios2_fast_data_master_byteenable                   (nios2_fast_data_master_byteenable),                        //                                              .byteenable
		.nios2_fast_data_master_read                         (nios2_fast_data_master_read),                              //                                              .read
		.nios2_fast_data_master_readdata                     (nios2_fast_data_master_readdata),                          //                                              .readdata
		.nios2_fast_data_master_readdatavalid                (nios2_fast_data_master_readdatavalid),                     //                                              .readdatavalid
		.nios2_fast_data_master_write                        (nios2_fast_data_master_write),                             //                                              .write
		.nios2_fast_data_master_writedata                    (nios2_fast_data_master_writedata),                         //                                              .writedata
		.nios2_fast_data_master_debugaccess                  (nios2_fast_data_master_debugaccess),                       //                                              .debugaccess
		.nios2_fast_instruction_master_address               (nios2_fast_instruction_master_address),                    //                 nios2_fast_instruction_master.address
		.nios2_fast_instruction_master_waitrequest           (nios2_fast_instruction_master_waitrequest),                //                                              .waitrequest
		.nios2_fast_instruction_master_read                  (nios2_fast_instruction_master_read),                       //                                              .read
		.nios2_fast_instruction_master_readdata              (nios2_fast_instruction_master_readdata),                   //                                              .readdata
		.nios2_fast_instruction_master_readdatavalid         (nios2_fast_instruction_master_readdatavalid),              //                                              .readdatavalid
		.peridot_hostbridge_m1_address                       (peridot_hostbridge_m1_address),                            //                         peridot_hostbridge_m1.address
		.peridot_hostbridge_m1_waitrequest                   (peridot_hostbridge_m1_waitrequest),                        //                                              .waitrequest
		.peridot_hostbridge_m1_byteenable                    (peridot_hostbridge_m1_byteenable),                         //                                              .byteenable
		.peridot_hostbridge_m1_read                          (peridot_hostbridge_m1_read),                               //                                              .read
		.peridot_hostbridge_m1_readdata                      (peridot_hostbridge_m1_readdata),                           //                                              .readdata
		.peridot_hostbridge_m1_readdatavalid                 (peridot_hostbridge_m1_readdatavalid),                      //                                              .readdatavalid
		.peridot_hostbridge_m1_write                         (peridot_hostbridge_m1_write),                              //                                              .write
		.peridot_hostbridge_m1_writedata                     (peridot_hostbridge_m1_writedata),                          //                                              .writedata
		.nios2_fast_debug_mem_slave_address                  (mm_interconnect_0_nios2_fast_debug_mem_slave_address),     //                    nios2_fast_debug_mem_slave.address
		.nios2_fast_debug_mem_slave_write                    (mm_interconnect_0_nios2_fast_debug_mem_slave_write),       //                                              .write
		.nios2_fast_debug_mem_slave_read                     (mm_interconnect_0_nios2_fast_debug_mem_slave_read),        //                                              .read
		.nios2_fast_debug_mem_slave_readdata                 (mm_interconnect_0_nios2_fast_debug_mem_slave_readdata),    //                                              .readdata
		.nios2_fast_debug_mem_slave_writedata                (mm_interconnect_0_nios2_fast_debug_mem_slave_writedata),   //                                              .writedata
		.nios2_fast_debug_mem_slave_byteenable               (mm_interconnect_0_nios2_fast_debug_mem_slave_byteenable),  //                                              .byteenable
		.nios2_fast_debug_mem_slave_waitrequest              (mm_interconnect_0_nios2_fast_debug_mem_slave_waitrequest), //                                              .waitrequest
		.nios2_fast_debug_mem_slave_debugaccess              (mm_interconnect_0_nios2_fast_debug_mem_slave_debugaccess), //                                              .debugaccess
		.peripheral_bridge_s0_address                        (mm_interconnect_0_peripheral_bridge_s0_address),           //                          peripheral_bridge_s0.address
		.peripheral_bridge_s0_write                          (mm_interconnect_0_peripheral_bridge_s0_write),             //                                              .write
		.peripheral_bridge_s0_read                           (mm_interconnect_0_peripheral_bridge_s0_read),              //                                              .read
		.peripheral_bridge_s0_readdata                       (mm_interconnect_0_peripheral_bridge_s0_readdata),          //                                              .readdata
		.peripheral_bridge_s0_writedata                      (mm_interconnect_0_peripheral_bridge_s0_writedata),         //                                              .writedata
		.peripheral_bridge_s0_burstcount                     (mm_interconnect_0_peripheral_bridge_s0_burstcount),        //                                              .burstcount
		.peripheral_bridge_s0_byteenable                     (mm_interconnect_0_peripheral_bridge_s0_byteenable),        //                                              .byteenable
		.peripheral_bridge_s0_readdatavalid                  (mm_interconnect_0_peripheral_bridge_s0_readdatavalid),     //                                              .readdatavalid
		.peripheral_bridge_s0_waitrequest                    (mm_interconnect_0_peripheral_bridge_s0_waitrequest),       //                                              .waitrequest
		.peripheral_bridge_s0_debugaccess                    (mm_interconnect_0_peripheral_bridge_s0_debugaccess),       //                                              .debugaccess
		.sdram_s1_address                                    (mm_interconnect_0_sdram_s1_address),                       //                                      sdram_s1.address
		.sdram_s1_write                                      (mm_interconnect_0_sdram_s1_write),                         //                                              .write
		.sdram_s1_read                                       (mm_interconnect_0_sdram_s1_read),                          //                                              .read
		.sdram_s1_readdata                                   (mm_interconnect_0_sdram_s1_readdata),                      //                                              .readdata
		.sdram_s1_writedata                                  (mm_interconnect_0_sdram_s1_writedata),                     //                                              .writedata
		.sdram_s1_byteenable                                 (mm_interconnect_0_sdram_s1_byteenable),                    //                                              .byteenable
		.sdram_s1_readdatavalid                              (mm_interconnect_0_sdram_s1_readdatavalid),                 //                                              .readdatavalid
		.sdram_s1_waitrequest                                (mm_interconnect_0_sdram_s1_waitrequest),                   //                                              .waitrequest
		.sdram_s1_chipselect                                 (mm_interconnect_0_sdram_s1_chipselect),                    //                                              .chipselect
		.ufm_data_address                                    (mm_interconnect_0_ufm_data_address),                       //                                      ufm_data.address
		.ufm_data_write                                      (mm_interconnect_0_ufm_data_write),                         //                                              .write
		.ufm_data_read                                       (mm_interconnect_0_ufm_data_read),                          //                                              .read
		.ufm_data_readdata                                   (mm_interconnect_0_ufm_data_readdata),                      //                                              .readdata
		.ufm_data_writedata                                  (mm_interconnect_0_ufm_data_writedata),                     //                                              .writedata
		.ufm_data_burstcount                                 (mm_interconnect_0_ufm_data_burstcount),                    //                                              .burstcount
		.ufm_data_readdatavalid                              (mm_interconnect_0_ufm_data_readdatavalid),                 //                                              .readdatavalid
		.ufm_data_waitrequest                                (mm_interconnect_0_ufm_data_waitrequest)                    //                                              .waitrequest
	);

	ngs_boot_core_mm_interconnect_1 mm_interconnect_1 (
		.core_clk_clk_clk                                    (clk_100m_clk),                                              //                                  core_clk_clk.clk
		.peri_clk_clk_clk                                    (clk_25m_clk),                                               //                                  peri_clk_clk.clk
		.jtag_uart_reset_reset_bridge_in_reset_reset         (rst_controller_001_reset_out_reset),                        //         jtag_uart_reset_reset_bridge_in_reset.reset
		.peripheral_bridge_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                            // peripheral_bridge_reset_reset_bridge_in_reset.reset
		.ufm_nreset_reset_bridge_in_reset_reset              (rst_controller_002_reset_out_reset),                        //              ufm_nreset_reset_bridge_in_reset.reset
		.peripheral_bridge_m0_address                        (peripheral_bridge_m0_address),                              //                          peripheral_bridge_m0.address
		.peripheral_bridge_m0_waitrequest                    (peripheral_bridge_m0_waitrequest),                          //                                              .waitrequest
		.peripheral_bridge_m0_burstcount                     (peripheral_bridge_m0_burstcount),                           //                                              .burstcount
		.peripheral_bridge_m0_byteenable                     (peripheral_bridge_m0_byteenable),                           //                                              .byteenable
		.peripheral_bridge_m0_read                           (peripheral_bridge_m0_read),                                 //                                              .read
		.peripheral_bridge_m0_readdata                       (peripheral_bridge_m0_readdata),                             //                                              .readdata
		.peripheral_bridge_m0_readdatavalid                  (peripheral_bridge_m0_readdatavalid),                        //                                              .readdatavalid
		.peripheral_bridge_m0_write                          (peripheral_bridge_m0_write),                                //                                              .write
		.peripheral_bridge_m0_writedata                      (peripheral_bridge_m0_writedata),                            //                                              .writedata
		.peripheral_bridge_m0_debugaccess                    (peripheral_bridge_m0_debugaccess),                          //                                              .debugaccess
		.gpio_s1_address                                     (mm_interconnect_1_gpio_s1_address),                         //                                       gpio_s1.address
		.gpio_s1_write                                       (mm_interconnect_1_gpio_s1_write),                           //                                              .write
		.gpio_s1_readdata                                    (mm_interconnect_1_gpio_s1_readdata),                        //                                              .readdata
		.gpio_s1_writedata                                   (mm_interconnect_1_gpio_s1_writedata),                       //                                              .writedata
		.gpio_s1_chipselect                                  (mm_interconnect_1_gpio_s1_chipselect),                      //                                              .chipselect
		.jtag_uart_avalon_jtag_slave_address                 (mm_interconnect_1_jtag_uart_avalon_jtag_slave_address),     //                   jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                   (mm_interconnect_1_jtag_uart_avalon_jtag_slave_write),       //                                              .write
		.jtag_uart_avalon_jtag_slave_read                    (mm_interconnect_1_jtag_uart_avalon_jtag_slave_read),        //                                              .read
		.jtag_uart_avalon_jtag_slave_readdata                (mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata),    //                                              .readdata
		.jtag_uart_avalon_jtag_slave_writedata               (mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata),   //                                              .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest             (mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest), //                                              .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect              (mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect),  //                                              .chipselect
		.peridot_hostbridge_s1_address                       (mm_interconnect_1_peridot_hostbridge_s1_address),           //                         peridot_hostbridge_s1.address
		.peridot_hostbridge_s1_write                         (mm_interconnect_1_peridot_hostbridge_s1_write),             //                                              .write
		.peridot_hostbridge_s1_read                          (mm_interconnect_1_peridot_hostbridge_s1_read),              //                                              .read
		.peridot_hostbridge_s1_readdata                      (mm_interconnect_1_peridot_hostbridge_s1_readdata),          //                                              .readdata
		.peridot_hostbridge_s1_writedata                     (mm_interconnect_1_peridot_hostbridge_s1_writedata),         //                                              .writedata
		.systimer_s1_address                                 (mm_interconnect_1_systimer_s1_address),                     //                                   systimer_s1.address
		.systimer_s1_write                                   (mm_interconnect_1_systimer_s1_write),                       //                                              .write
		.systimer_s1_readdata                                (mm_interconnect_1_systimer_s1_readdata),                    //                                              .readdata
		.systimer_s1_writedata                               (mm_interconnect_1_systimer_s1_writedata),                   //                                              .writedata
		.systimer_s1_chipselect                              (mm_interconnect_1_systimer_s1_chipselect),                  //                                              .chipselect
		.ufm_csr_address                                     (mm_interconnect_1_ufm_csr_address),                         //                                       ufm_csr.address
		.ufm_csr_write                                       (mm_interconnect_1_ufm_csr_write),                           //                                              .write
		.ufm_csr_read                                        (mm_interconnect_1_ufm_csr_read),                            //                                              .read
		.ufm_csr_readdata                                    (mm_interconnect_1_ufm_csr_readdata),                        //                                              .readdata
		.ufm_csr_writedata                                   (mm_interconnect_1_ufm_csr_writedata)                        //                                              .writedata
	);

	ngs_boot_core_irq_mapper irq_mapper (
		.clk           (clk_100m_clk),                       //       clk.clk
		.reset         (rst_controller_002_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.sender_irq    (nios2_fast_irq_irq)                  //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (clk_25m_clk),                        //       receiver_clk.clk
		.sender_clk     (clk_100m_clk),                       //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_002_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver1_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_001 (
		.receiver_clk   (clk_25m_clk),                        //       receiver_clk.clk
		.sender_clk     (clk_100m_clk),                       //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_002_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_001_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver3_irq)            //             sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_25m_clk),                    //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_100m_clk),                       //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.clk            (clk_100m_clk),                           //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_002_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
